module InitialPermutation(input [63:0] dataIn, output [63:0] dataOut);
    assign dataOut[ 0] = dataIn[57];
    assign dataOut[ 1] = dataIn[49];
    assign dataOut[ 2] = dataIn[41];
    assign dataOut[ 3] = dataIn[33];
    assign dataOut[ 4] = dataIn[25];
    assign dataOut[ 5] = dataIn[17];
    assign dataOut[ 6] = dataIn[ 9];
    assign dataOut[ 7] = dataIn[ 1];
    assign dataOut[ 8] = dataIn[59];
    assign dataOut[ 9] = dataIn[51];
    assign dataOut[10] = dataIn[43];
    assign dataOut[11] = dataIn[35];
    assign dataOut[12] = dataIn[27];
    assign dataOut[13] = dataIn[19];
    assign dataOut[14] = dataIn[11];
    assign dataOut[15] = dataIn[ 3];
    assign dataOut[16] = dataIn[61];
    assign dataOut[17] = dataIn[53];
    assign dataOut[18] = dataIn[45];
    assign dataOut[19] = dataIn[37];
    assign dataOut[20] = dataIn[29];
    assign dataOut[21] = dataIn[21];
    assign dataOut[22] = dataIn[13];
    assign dataOut[23] = dataIn[ 5];
    assign dataOut[24] = dataIn[63];
    assign dataOut[25] = dataIn[55];
    assign dataOut[26] = dataIn[47];
    assign dataOut[27] = dataIn[39];
    assign dataOut[28] = dataIn[31];
    assign dataOut[29] = dataIn[23];
    assign dataOut[30] = dataIn[15];
    assign dataOut[31] = dataIn[ 7];
    assign dataOut[32] = dataIn[56];
    assign dataOut[33] = dataIn[48];
    assign dataOut[34] = dataIn[40];
    assign dataOut[35] = dataIn[32];
    assign dataOut[36] = dataIn[24];
    assign dataOut[37] = dataIn[16];
    assign dataOut[38] = dataIn[ 8];
    assign dataOut[39] = dataIn[ 0];
    assign dataOut[40] = dataIn[58];
    assign dataOut[41] = dataIn[50];
    assign dataOut[42] = dataIn[42];
    assign dataOut[43] = dataIn[34];
    assign dataOut[44] = dataIn[26];
    assign dataOut[45] = dataIn[18];
    assign dataOut[46] = dataIn[10];
    assign dataOut[47] = dataIn[ 2];
    assign dataOut[48] = dataIn[60];
    assign dataOut[49] = dataIn[52];
    assign dataOut[50] = dataIn[44];
    assign dataOut[51] = dataIn[36];
    assign dataOut[52] = dataIn[28];
    assign dataOut[53] = dataIn[20];
    assign dataOut[54] = dataIn[12];
    assign dataOut[55] = dataIn[ 4];
    assign dataOut[56] = dataIn[62];
    assign dataOut[57] = dataIn[54];
    assign dataOut[58] = dataIn[46];
    assign dataOut[59] = dataIn[38];
    assign dataOut[60] = dataIn[30];
    assign dataOut[61] = dataIn[22];
    assign dataOut[62] = dataIn[14];
    assign dataOut[63] = dataIn[ 6];
endmodule
module FinalPermutation(input [63:0] dataIn, output [63:0] dataOut);
    assign dataOut[ 0] = dataIn[39];
    assign dataOut[ 1] = dataIn[ 7];
    assign dataOut[ 2] = dataIn[47];
    assign dataOut[ 3] = dataIn[15];
    assign dataOut[ 4] = dataIn[55];
    assign dataOut[ 5] = dataIn[23];
    assign dataOut[ 6] = dataIn[63];
    assign dataOut[ 7] = dataIn[31];
    assign dataOut[ 8] = dataIn[38];
    assign dataOut[ 9] = dataIn[ 6];
    assign dataOut[10] = dataIn[46];
    assign dataOut[11] = dataIn[14];
    assign dataOut[12] = dataIn[54];
    assign dataOut[13] = dataIn[22];
    assign dataOut[14] = dataIn[62];
    assign dataOut[15] = dataIn[30];
    assign dataOut[16] = dataIn[37];
    assign dataOut[17] = dataIn[ 5];
    assign dataOut[18] = dataIn[45];
    assign dataOut[19] = dataIn[13];
    assign dataOut[20] = dataIn[53];
    assign dataOut[21] = dataIn[21];
    assign dataOut[22] = dataIn[61];
    assign dataOut[23] = dataIn[29];
    assign dataOut[24] = dataIn[36];
    assign dataOut[25] = dataIn[ 4];
    assign dataOut[26] = dataIn[44];
    assign dataOut[27] = dataIn[12];
    assign dataOut[28] = dataIn[52];
    assign dataOut[29] = dataIn[20];
    assign dataOut[30] = dataIn[60];
    assign dataOut[31] = dataIn[28];
    assign dataOut[32] = dataIn[35];
    assign dataOut[33] = dataIn[ 3];
    assign dataOut[34] = dataIn[43];
    assign dataOut[35] = dataIn[11];
    assign dataOut[36] = dataIn[51];
    assign dataOut[37] = dataIn[19];
    assign dataOut[38] = dataIn[59];
    assign dataOut[39] = dataIn[27];
    assign dataOut[40] = dataIn[34];
    assign dataOut[41] = dataIn[ 2];
    assign dataOut[42] = dataIn[42];
    assign dataOut[43] = dataIn[10];
    assign dataOut[44] = dataIn[50];
    assign dataOut[45] = dataIn[18];
    assign dataOut[46] = dataIn[58];
    assign dataOut[47] = dataIn[26];
    assign dataOut[48] = dataIn[33];
    assign dataOut[49] = dataIn[ 1];
    assign dataOut[50] = dataIn[41];
    assign dataOut[51] = dataIn[ 9];
    assign dataOut[52] = dataIn[49];
    assign dataOut[53] = dataIn[17];
    assign dataOut[54] = dataIn[57];
    assign dataOut[55] = dataIn[25];
    assign dataOut[56] = dataIn[32];
    assign dataOut[57] = dataIn[ 0];
    assign dataOut[58] = dataIn[40];
    assign dataOut[59] = dataIn[ 8];
    assign dataOut[60] = dataIn[48];
    assign dataOut[61] = dataIn[16];
    assign dataOut[62] = dataIn[56];
    assign dataOut[63] = dataIn[24];
endmodule
module ExpansionDBoxTable(input [31:0] dataIn, output [47:0] dataOut);
    assign dataOut[ 0] = dataIn[31];
    assign dataOut[ 1] = dataIn[ 0];
    assign dataOut[ 2] = dataIn[ 1];
    assign dataOut[ 3] = dataIn[ 2];
    assign dataOut[ 4] = dataIn[ 3];
    assign dataOut[ 5] = dataIn[ 4];
    assign dataOut[ 6] = dataIn[ 3];
    assign dataOut[ 7] = dataIn[ 4];
    assign dataOut[ 8] = dataIn[ 5];
    assign dataOut[ 9] = dataIn[ 6];
    assign dataOut[10] = dataIn[ 7];
    assign dataOut[11] = dataIn[ 8];
    assign dataOut[12] = dataIn[ 7];
    assign dataOut[13] = dataIn[ 8];
    assign dataOut[14] = dataIn[ 9];
    assign dataOut[15] = dataIn[10];
    assign dataOut[16] = dataIn[11];
    assign dataOut[17] = dataIn[12];
    assign dataOut[18] = dataIn[11];
    assign dataOut[19] = dataIn[12];
    assign dataOut[20] = dataIn[13];
    assign dataOut[21] = dataIn[14];
    assign dataOut[22] = dataIn[15];
    assign dataOut[23] = dataIn[16];
    assign dataOut[24] = dataIn[15];
    assign dataOut[25] = dataIn[16];
    assign dataOut[26] = dataIn[17];
    assign dataOut[27] = dataIn[18];
    assign dataOut[28] = dataIn[19];
    assign dataOut[29] = dataIn[20];
    assign dataOut[30] = dataIn[19];
    assign dataOut[31] = dataIn[20];
    assign dataOut[32] = dataIn[21];
    assign dataOut[33] = dataIn[22];
    assign dataOut[34] = dataIn[23];
    assign dataOut[35] = dataIn[24];
    assign dataOut[36] = dataIn[23];
    assign dataOut[37] = dataIn[24];
    assign dataOut[38] = dataIn[25];
    assign dataOut[39] = dataIn[26];
    assign dataOut[40] = dataIn[27];
    assign dataOut[41] = dataIn[28];
    assign dataOut[42] = dataIn[27];
    assign dataOut[43] = dataIn[28];
    assign dataOut[44] = dataIn[30];
    assign dataOut[45] = dataIn[30];
    assign dataOut[46] = dataIn[31];
    assign dataOut[47] = dataIn[ 0];
endmodule
module StraightDBoxTable(input [31:0] dataIn, output [31:0] dataOut);
    assign dataOut[ 0] = dataIn[15];
    assign dataOut[ 1] = dataIn[ 6];
    assign dataOut[ 2] = dataIn[19];
    assign dataOut[ 3] = dataIn[20];
    assign dataOut[ 4] = dataIn[28];
    assign dataOut[ 5] = dataIn[11];
    assign dataOut[ 6] = dataIn[27];
    assign dataOut[ 7] = dataIn[16];
    assign dataOut[ 8] = dataIn[ 0];
    assign dataOut[ 9] = dataIn[14];
    assign dataOut[10] = dataIn[22];
    assign dataOut[11] = dataIn[25];
    assign dataOut[12] = dataIn[ 4];
    assign dataOut[13] = dataIn[17];
    assign dataOut[14] = dataIn[30];
    assign dataOut[15] = dataIn[ 9];
    assign dataOut[16] = dataIn[ 1];
    assign dataOut[17] = dataIn[ 7];
    assign dataOut[18] = dataIn[23];
    assign dataOut[19] = dataIn[13];
    assign dataOut[20] = dataIn[31];
    assign dataOut[21] = dataIn[26];
    assign dataOut[22] = dataIn[ 2];
    assign dataOut[23] = dataIn[ 8];
    assign dataOut[24] = dataIn[18];
    assign dataOut[25] = dataIn[12];
    assign dataOut[26] = dataIn[29];
    assign dataOut[27] = dataIn[ 5];
    assign dataOut[28] = dataIn[21];
    assign dataOut[29] = dataIn[10];
    assign dataOut[30] = dataIn[ 3];
    assign dataOut[31] = dataIn[24];
endmodule
module ParityBitDropTable(input [63:0] dataIn, output [55:0] dataOut);
    assign dataOut[ 0] = dataIn[56];
    assign dataOut[ 1] = dataIn[48];
    assign dataOut[ 2] = dataIn[40];
    assign dataOut[ 3] = dataIn[32];
    assign dataOut[ 4] = dataIn[24];
    assign dataOut[ 5] = dataIn[16];
    assign dataOut[ 6] = dataIn[ 8];
    assign dataOut[ 7] = dataIn[ 0];
    assign dataOut[ 8] = dataIn[57];
    assign dataOut[ 9] = dataIn[49];
    assign dataOut[10] = dataIn[41];
    assign dataOut[11] = dataIn[33];
    assign dataOut[12] = dataIn[25];
    assign dataOut[13] = dataIn[17];
    assign dataOut[14] = dataIn[ 9];
    assign dataOut[15] = dataIn[ 1];
    assign dataOut[16] = dataIn[58];
    assign dataOut[17] = dataIn[50];
    assign dataOut[18] = dataIn[42];
    assign dataOut[19] = dataIn[34];
    assign dataOut[20] = dataIn[26];
    assign dataOut[21] = dataIn[18];
    assign dataOut[22] = dataIn[10];
    assign dataOut[23] = dataIn[ 2];
    assign dataOut[24] = dataIn[59];
    assign dataOut[25] = dataIn[51];
    assign dataOut[26] = dataIn[43];
    assign dataOut[27] = dataIn[35];
    assign dataOut[28] = dataIn[62];
    assign dataOut[29] = dataIn[54];
    assign dataOut[30] = dataIn[46];
    assign dataOut[31] = dataIn[38];
    assign dataOut[32] = dataIn[30];
    assign dataOut[33] = dataIn[22];
    assign dataOut[34] = dataIn[14];
    assign dataOut[35] = dataIn[ 6];
    assign dataOut[36] = dataIn[61];
    assign dataOut[37] = dataIn[53];
    assign dataOut[38] = dataIn[45];
    assign dataOut[39] = dataIn[37];
    assign dataOut[40] = dataIn[29];
    assign dataOut[41] = dataIn[21];
    assign dataOut[42] = dataIn[13];
    assign dataOut[43] = dataIn[ 5];
    assign dataOut[44] = dataIn[60];
    assign dataOut[45] = dataIn[52];
    assign dataOut[46] = dataIn[44];
    assign dataOut[47] = dataIn[36];
    assign dataOut[48] = dataIn[28];
    assign dataOut[49] = dataIn[20];
    assign dataOut[50] = dataIn[12];
    assign dataOut[51] = dataIn[ 4];
    assign dataOut[52] = dataIn[27];
    assign dataOut[53] = dataIn[19];
    assign dataOut[54] = dataIn[11];
    assign dataOut[55] = dataIn[ 3];
endmodule
module KeyCompressionTable(input [55:0] dataIn, output [47:0] dataOut);
    assign dataOut[ 0] = dataIn[13];
    assign dataOut[ 1] = dataIn[16];
    assign dataOut[ 2] = dataIn[10];
    assign dataOut[ 3] = dataIn[23];
    assign dataOut[ 4] = dataIn[ 0];
    assign dataOut[ 5] = dataIn[ 4];
    assign dataOut[ 6] = dataIn[ 2];
    assign dataOut[ 7] = dataIn[27];
    assign dataOut[ 8] = dataIn[14];
    assign dataOut[ 9] = dataIn[ 5];
    assign dataOut[10] = dataIn[20];
    assign dataOut[11] = dataIn[ 9];
    assign dataOut[12] = dataIn[22];
    assign dataOut[13] = dataIn[18];
    assign dataOut[14] = dataIn[11];
    assign dataOut[15] = dataIn[ 3];
    assign dataOut[16] = dataIn[25];
    assign dataOut[17] = dataIn[ 7];
    assign dataOut[18] = dataIn[15];
    assign dataOut[19] = dataIn[ 6];
    assign dataOut[20] = dataIn[26];
    assign dataOut[21] = dataIn[19];
    assign dataOut[22] = dataIn[12];
    assign dataOut[23] = dataIn[ 1];
    assign dataOut[24] = dataIn[40];
    assign dataOut[25] = dataIn[51];
    assign dataOut[26] = dataIn[30];
    assign dataOut[27] = dataIn[36];
    assign dataOut[28] = dataIn[46];
    assign dataOut[29] = dataIn[54];
    assign dataOut[30] = dataIn[29];
    assign dataOut[31] = dataIn[39];
    assign dataOut[32] = dataIn[50];
    assign dataOut[33] = dataIn[44];
    assign dataOut[34] = dataIn[32];
    assign dataOut[35] = dataIn[47];
    assign dataOut[36] = dataIn[43];
    assign dataOut[37] = dataIn[48];
    assign dataOut[38] = dataIn[38];
    assign dataOut[39] = dataIn[55];
    assign dataOut[40] = dataIn[33];
    assign dataOut[41] = dataIn[52];
    assign dataOut[42] = dataIn[45];
    assign dataOut[43] = dataIn[41];
    assign dataOut[44] = dataIn[49];
    assign dataOut[45] = dataIn[35];
    assign dataOut[46] = dataIn[28];
    assign dataOut[47] = dataIn[31];
endmodule
